module and16 (
    input [15:0] a,
    output y
);
    assign y = &a;
endmodule